module rx_fsm(
    input logic clk, nRST,
    
);